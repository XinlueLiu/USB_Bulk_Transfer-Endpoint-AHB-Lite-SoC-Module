module flex_pts_sr
#(
parameter NUM_BITS = 4,
parameter SHIFT_MSB = 1
)
(
input wire clk,
input wire n_rst,
input wire shift_enable,
input wire load_enable,
input wire halt,
input wire[NUM_BITS-1:0] parallel_in,
output reg serial_out,
output reg [NUM_BITS-1:0]parallel_out
);
integer i;
reg new_serial_out;
reg [NUM_BITS-1:0] new_parallel_out;
//reg [NUM_BITS:0] parallel_out;
always_ff @(posedge clk,negedge n_rst)
begin 
	if(n_rst == 1'b0) begin
		serial_out <= '0;
	end
	else begin
		serial_out <=new_serial_out;
		parallel_out<=new_parallel_out;
	end
end
always_comb
begin
   if(halt == 1'b1) begin
	new_serial_out = serial_out;
	new_parallel_out = parallel_out;
   end
  else begin
   if(load_enable == 1'b1)
    	begin
	new_parallel_out[NUM_BITS-2:0] = parallel_in[NUM_BITS-1:1];
	new_serial_out = parallel_in[0];
	new_parallel_out[NUM_BITS-1] = 0;
	end
  	 else begin
		if(shift_enable == 1'b1)
		begin
 	  		if(SHIFT_MSB == 1)
	 		 begin
	 		new_parallel_out[0] = 0;
			/*for(i = 1;i<=NUM_BITS-1 ; i = i+1)
			begin
			new_parallel_out[i] = parallel_out[i-1];
			end*/
			new_parallel_out[NUM_BITS-1:1] = parallel_out[NUM_BITS-2:0];
			new_parallel_out[0] = 0;
			new_serial_out = new_parallel_out[NUM_BITS-1];
 	  		end
	  		else begin

			new_parallel_out[NUM_BITS-1] = 0;
			/*for(i = 0;i<=NUM_BITS-2 ; i = i+1)
			begin
			new_parallel_out[i] = parallel_out[i+1];
			end*/
			//endgenerate
			new_parallel_out[NUM_BITS-2:0] = parallel_out[NUM_BITS-1:1];
			new_serial_out = parallel_out[0];
	   		end
	  	end
		else begin
			new_parallel_out = parallel_out;
			new_serial_out = serial_out;
		end
	end
   end
end
endmodule
